module Processor(input_dummy, output_dummy);
input input_dummy;
output output_dummy;

assign output_dummy = !input_dummy;
endmodule